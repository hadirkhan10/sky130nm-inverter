magic
tech sky130A
timestamp 1647808945
<< nwell >>
rect -56 -48 107 98
<< nmos >>
rect 34 -140 49 -98
<< pmos >>
rect 34 -30 49 54
<< ndiff >>
rect -2 -115 34 -98
rect -2 -132 2 -115
rect 19 -132 34 -115
rect -2 -140 34 -132
rect 49 -106 85 -98
rect 49 -123 64 -106
rect 81 -123 85 -106
rect 49 -140 85 -123
<< pdiff >>
rect 4 34 34 54
rect 4 1 8 34
rect 25 1 34 34
rect 4 -30 34 1
rect 49 34 83 54
rect 49 1 62 34
rect 79 1 83 34
rect 49 -30 83 1
<< ndiffc >>
rect 2 -132 19 -115
rect 64 -123 81 -106
<< pdiffc >>
rect 8 1 25 34
rect 62 1 79 34
<< psubdiff >>
rect -37 -111 -2 -98
rect -37 -128 -32 -111
rect -15 -128 -2 -111
rect -37 -140 -2 -128
<< nsubdiff >>
rect -38 32 4 54
rect -38 -1 -26 32
rect -9 -1 4 32
rect -38 -30 4 -1
<< psubdiffcont >>
rect -32 -128 -15 -111
<< nsubdiffcont >>
rect -26 -1 -9 32
<< poly >>
rect 34 54 49 67
rect 34 -52 49 -30
rect 0 -57 49 -52
rect 0 -74 8 -57
rect 26 -74 49 -57
rect 0 -79 49 -74
rect 34 -98 49 -79
rect 34 -165 49 -140
<< polycont >>
rect 8 -74 26 -57
<< locali >>
rect 4 94 25 95
rect 4 77 6 94
rect 23 77 25 94
rect 4 40 25 77
rect -28 34 25 40
rect -28 32 8 34
rect -28 -1 -26 32
rect -9 1 8 32
rect -9 -1 25 1
rect -28 -10 25 -1
rect 4 -30 25 -10
rect 62 34 83 54
rect 79 1 83 34
rect 62 -30 83 1
rect 0 -57 34 -52
rect 0 -74 8 -57
rect 26 -74 34 -57
rect 0 -79 34 -74
rect 64 -53 83 -30
rect 64 -58 117 -53
rect 64 -75 91 -58
rect 109 -75 117 -58
rect 64 -80 117 -75
rect 64 -98 83 -80
rect -37 -111 21 -103
rect -37 -128 -32 -111
rect -15 -115 21 -111
rect -15 -128 2 -115
rect -37 -132 2 -128
rect 19 -132 21 -115
rect -37 -140 21 -132
rect 62 -106 85 -98
rect 62 -123 64 -106
rect 81 -123 85 -106
rect 62 -140 85 -123
rect -2 -157 21 -140
rect -2 -174 1 -157
rect 18 -174 21 -157
rect -2 -176 21 -174
<< viali >>
rect 6 77 23 94
rect 8 -74 26 -57
rect 91 -75 109 -58
rect 1 -174 18 -157
<< metal1 >>
rect -61 94 112 98
rect -61 77 6 94
rect 23 77 112 94
rect -61 74 112 77
rect 0 -57 34 -52
rect 0 -74 8 -57
rect 26 -74 34 -57
rect 0 -79 34 -74
rect 83 -58 117 -53
rect 83 -75 91 -58
rect 109 -75 117 -58
rect 83 -80 117 -75
rect -61 -157 112 -154
rect -61 -174 1 -157
rect 18 -174 112 -157
rect -61 -178 112 -174
<< labels >>
rlabel metal1 15 -70 21 -63 1 A
port 1 n
rlabel viali 97 -70 104 -63 1 Z
port 2 n
rlabel viali 12 84 16 88 1 VDD
port 5 n
rlabel viali 7 -168 12 -162 1 GND
port 6 n
<< end >>
