* NGSPICE file created from INV.ext - technology: sky130A

.subckt INV A Z VDD GND
X0 Z A VDD VDD sky130_fd_pr__pfet_01v8 ad=2.856e+11p pd=2.36e+06u as=2.52e+11p ps=2.28e+06u w=840000u l=150000u
X1 Z A GND GND sky130_fd_pr__nfet_01v8 ad=1.512e+11p pd=1.56e+06u as=1.512e+11p ps=1.56e+06u w=420000u l=150000u
.ends

